    0  => x"20030001",
    1  => x"00032820",
    2  => x"00a33822",
    3  => x"20640004",
    4  => x"00641024",
    5  => x"00472825",
    6  => x"10e30008",
    7  => x"00000020",
    8  => x"00000020",
    9  => x"0085102a",
    10  => x"ac841fd7",
    11  => x"8ca21fdb",
    12  => x"2047fffc",
    13  => x"08000006",
    14  => x"00000020",
    15  => x"00e2202a",
    16  => x"00e31024",
    17  => x"8c471fdb",
    18  => x"ac452003",
    19  => x"10a70003",
    20  => x"00000020",
    21  => x"00000020",
    22  => x"00a33825",
    23  => x"8ce42003",
    24  => x"08000000",
    25  => x"00000020",
    26  => x"00000020",
